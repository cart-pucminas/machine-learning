ShiftReg_inst : ShiftReg PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		shiftout	 => shiftout_sig
	);
