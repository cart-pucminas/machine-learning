Kmeans_RomMemory_inst : Kmeans_RomMemory PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
