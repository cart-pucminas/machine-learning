-- megafunction wizard: %ALTFP_COMPARE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_compare 

-- ============================================================
-- File Name: CompareALessB.vhd
-- Megafunction Name(s):
-- 			altfp_compare
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_compare CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone III" PIPELINE=1 WIDTH_EXP=8 WIDTH_MAN=23 alb clk_en clock dataa datab
--VERSION_BEGIN 9.1SP2 cbx_altfp_compare 2010:03:24:20:43:42:SJ cbx_cycloneii 2010:03:24:20:43:43:SJ cbx_lpm_add_sub 2010:03:24:20:43:43:SJ cbx_lpm_compare 2010:03:24:20:43:43:SJ cbx_mgl 2010:03:24:21:01:05:SJ cbx_stratix 2010:03:24:20:43:43:SJ cbx_stratixii 2010:03:24:20:43:43:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 4 reg 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  CompareALessB_altfp_compare_ksb IS 
	 PORT 
	 ( 
		 alb	:	OUT  STD_LOGIC;
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END CompareALessB_altfp_compare_ksb;

 ARCHITECTURE RTL OF CompareALessB_altfp_compare_ksb IS

	 SIGNAL	 out_alb_w_dffe3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cmpr1_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr1_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr2_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr2_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_agb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w304w305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_agb_w_dffe2_wo314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_flip_outputs_dffe2_wo310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range11w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range21w28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range31w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range41w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range51w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range61w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range71w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range14w20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range24w30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range34w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range44w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range54w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range64w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range74w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_aeb_range233w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_aeb_range237w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_aeb_range241w250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range251w254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range251w260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range253w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range253w262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_eq_grp_range255w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_both_inputs_zero_dffe2_wo312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_a_not_zero_dffe1_wo293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_agb_w_dffe2_wo309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_b_not_zero_dffe1_wo294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_dataa_zero_w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_datab_zero_w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_out_aeb_w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_out_agb_w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_out_unordered_w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w304w305w306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range141w143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range147w149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range157w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range163w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range169w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range175w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range181w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range187w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range193w195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range87w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range199w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range205w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range211w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range11w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range21w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range31w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range41w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range51w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range61w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range93w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range71w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range99w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range105w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range111w113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range117w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range123w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range129w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range135w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range144w146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range150w152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range160w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range166w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range172w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range178w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range184w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range190w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range196w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range90w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range202w204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range208w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range214w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range14w16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range24w26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range34w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range44w46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range54w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range64w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range96w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range74w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range102w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range108w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range114w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range120w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range126w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range132w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range138w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_agb_tmp_w_range265w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_agb_tmp_w_range267w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_agb_tmp_w_range269w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_not_zero_dffe1_wo_range285w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_not_zero_dffe1_wo_range288w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_adjusted_dffe2_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_adjusted_dffe2_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_adjusted_w :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe1_wi :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_dffe1_wo :	STD_LOGIC;
	 SIGNAL  aligned_dataa_sign_w :	STD_LOGIC;
	 SIGNAL  aligned_dataa_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  aligned_datab_sign_adjusted_dffe2_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_adjusted_dffe2_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_adjusted_w :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe1_wi :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_dffe1_wo :	STD_LOGIC;
	 SIGNAL  aligned_datab_sign_w :	STD_LOGIC;
	 SIGNAL  aligned_datab_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  both_inputs_zero :	STD_LOGIC;
	 SIGNAL  both_inputs_zero_dffe2_wi :	STD_LOGIC;
	 SIGNAL  both_inputs_zero_dffe2_wo :	STD_LOGIC;
	 SIGNAL  exp_a_all_one_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_a_all_one_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_a_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_not_zero_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_a_not_zero_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_a_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_aeb :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_aeb_tmp_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_aeb_w :	STD_LOGIC;
	 SIGNAL  exp_aeb_w_dffe2_wi :	STD_LOGIC;
	 SIGNAL  exp_aeb_w_dffe2_wo :	STD_LOGIC;
	 SIGNAL  exp_agb :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_agb_tmp_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  exp_agb_w :	STD_LOGIC;
	 SIGNAL  exp_agb_w_dffe2_wi :	STD_LOGIC;
	 SIGNAL  exp_agb_w_dffe2_wo :	STD_LOGIC;
	 SIGNAL  exp_b_all_one_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_b_all_one_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_b_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_not_zero_dffe1_wi :	STD_LOGIC;
	 SIGNAL  exp_b_not_zero_dffe1_wo :	STD_LOGIC;
	 SIGNAL  exp_b_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_eq_grp :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  exp_eq_gt_grp :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  flip_outputs_dffe2_wi :	STD_LOGIC;
	 SIGNAL  flip_outputs_dffe2_wo :	STD_LOGIC;
	 SIGNAL  flip_outputs_w :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe2_wi :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_dffe2_wo :	STD_LOGIC;
	 SIGNAL  input_dataa_nan_w :	STD_LOGIC;
	 SIGNAL  input_dataa_zero_w :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe2_wi :	STD_LOGIC;
	 SIGNAL  input_datab_nan_dffe2_wo :	STD_LOGIC;
	 SIGNAL  input_datab_nan_w :	STD_LOGIC;
	 SIGNAL  input_datab_zero_w :	STD_LOGIC;
	 SIGNAL  man_a_not_zero_dffe1_wi :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_a_not_zero_dffe1_wo :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_a_not_zero_merge_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_a_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_not_zero_dffe1_wi :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_b_not_zero_dffe1_wo :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_b_not_zero_merge_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  man_b_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  out_aeb_w :	STD_LOGIC;
	 SIGNAL  out_agb_w :	STD_LOGIC;
	 SIGNAL  out_alb_dffe3_wi :	STD_LOGIC;
	 SIGNAL  out_alb_dffe3_wo :	STD_LOGIC;
	 SIGNAL  out_alb_w :	STD_LOGIC;
	 SIGNAL  out_unordered_w :	STD_LOGIC;
	 SIGNAL  wire_w_dataa_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_all_one_w_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_not_zero_w_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_range237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_tmp_w_range243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_tmp_w_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_aeb_tmp_w_range247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_range234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_range238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_tmp_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_tmp_w_range267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_agb_tmp_w_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_all_one_w_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_not_zero_w_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_grp_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_grp_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_grp_range255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_gt_grp_range259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_gt_grp_range261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_eq_gt_grp_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_dffe1_wo_range285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_merge_w_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_not_zero_w_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_dffe1_wo_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_merge_w_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_not_zero_w_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w304w305w(0) <= wire_w304w(0) AND exp_aeb_w_dffe2_wo;
	wire_w316w(0) <= wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w(0) AND aligned_datab_sign_adjusted_dffe2_wo;
	wire_w_lg_exp_agb_w_dffe2_wo314w(0) <= exp_agb_w_dffe2_wo AND wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w(0);
	wire_w_lg_flip_outputs_dffe2_wo310w(0) <= flip_outputs_dffe2_wo AND wire_w_lg_exp_agb_w_dffe2_wo309w(0);
	wire_w_lg_w_dataa_range11w18w(0) <= wire_w_dataa_range11w(0) AND wire_w_exp_a_all_one_w_range7w(0);
	wire_w_lg_w_dataa_range21w28w(0) <= wire_w_dataa_range21w(0) AND wire_w_exp_a_all_one_w_range17w(0);
	wire_w_lg_w_dataa_range31w38w(0) <= wire_w_dataa_range31w(0) AND wire_w_exp_a_all_one_w_range27w(0);
	wire_w_lg_w_dataa_range41w48w(0) <= wire_w_dataa_range41w(0) AND wire_w_exp_a_all_one_w_range37w(0);
	wire_w_lg_w_dataa_range51w58w(0) <= wire_w_dataa_range51w(0) AND wire_w_exp_a_all_one_w_range47w(0);
	wire_w_lg_w_dataa_range61w68w(0) <= wire_w_dataa_range61w(0) AND wire_w_exp_a_all_one_w_range57w(0);
	wire_w_lg_w_dataa_range71w78w(0) <= wire_w_dataa_range71w(0) AND wire_w_exp_a_all_one_w_range67w(0);
	wire_w_lg_w_datab_range14w20w(0) <= wire_w_datab_range14w(0) AND wire_w_exp_b_all_one_w_range9w(0);
	wire_w_lg_w_datab_range24w30w(0) <= wire_w_datab_range24w(0) AND wire_w_exp_b_all_one_w_range19w(0);
	wire_w_lg_w_datab_range34w40w(0) <= wire_w_datab_range34w(0) AND wire_w_exp_b_all_one_w_range29w(0);
	wire_w_lg_w_datab_range44w50w(0) <= wire_w_datab_range44w(0) AND wire_w_exp_b_all_one_w_range39w(0);
	wire_w_lg_w_datab_range54w60w(0) <= wire_w_datab_range54w(0) AND wire_w_exp_b_all_one_w_range49w(0);
	wire_w_lg_w_datab_range64w70w(0) <= wire_w_datab_range64w(0) AND wire_w_exp_b_all_one_w_range59w(0);
	wire_w_lg_w_datab_range74w80w(0) <= wire_w_datab_range74w(0) AND wire_w_exp_b_all_one_w_range69w(0);
	wire_w_lg_w_exp_aeb_range233w246w(0) <= wire_w_exp_aeb_range233w(0) AND wire_w_exp_aeb_tmp_w_range243w(0);
	wire_w_lg_w_exp_aeb_range237w248w(0) <= wire_w_exp_aeb_range237w(0) AND wire_w_exp_aeb_tmp_w_range245w(0);
	wire_w_lg_w_exp_aeb_range241w250w(0) <= wire_w_exp_aeb_range241w(0) AND wire_w_exp_aeb_tmp_w_range247w(0);
	wire_w_lg_w_exp_eq_grp_range251w254w(0) <= wire_w_exp_eq_grp_range251w(0) AND wire_w_exp_aeb_range233w(0);
	wire_w_lg_w_exp_eq_grp_range251w260w(0) <= wire_w_exp_eq_grp_range251w(0) AND wire_w_exp_agb_range234w(0);
	wire_w_lg_w_exp_eq_grp_range253w256w(0) <= wire_w_exp_eq_grp_range253w(0) AND wire_w_exp_aeb_range237w(0);
	wire_w_lg_w_exp_eq_grp_range253w262w(0) <= wire_w_exp_eq_grp_range253w(0) AND wire_w_exp_agb_range238w(0);
	wire_w_lg_w_exp_eq_grp_range255w264w(0) <= wire_w_exp_eq_grp_range255w(0) AND wire_w_exp_agb_range242w(0);
	wire_w304w(0) <= NOT wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo303w(0);
	wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo313w(0) <= NOT aligned_dataa_sign_adjusted_dffe2_wo;
	wire_w_lg_both_inputs_zero_dffe2_wo312w(0) <= NOT both_inputs_zero_dffe2_wo;
	wire_w_lg_exp_a_not_zero_dffe1_wo293w(0) <= NOT exp_a_not_zero_dffe1_wo;
	wire_w_lg_exp_agb_w_dffe2_wo309w(0) <= NOT exp_agb_w_dffe2_wo;
	wire_w_lg_exp_b_not_zero_dffe1_wo294w(0) <= NOT exp_b_not_zero_dffe1_wo;
	wire_w_lg_input_dataa_zero_w296w(0) <= NOT input_dataa_zero_w;
	wire_w_lg_input_datab_zero_w298w(0) <= NOT input_datab_zero_w;
	wire_w_lg_out_aeb_w308w(0) <= NOT out_aeb_w;
	wire_w_lg_out_agb_w320w(0) <= NOT out_agb_w;
	wire_w_lg_out_unordered_w302w(0) <= NOT out_unordered_w;
	wire_w_lg_w_lg_w304w305w306w(0) <= wire_w_lg_w304w305w(0) OR both_inputs_zero_dffe2_wo;
	wire_w_lg_w_dataa_range141w143w(0) <= wire_w_dataa_range141w(0) OR wire_w_man_a_not_zero_w_range136w(0);
	wire_w_lg_w_dataa_range147w149w(0) <= wire_w_dataa_range147w(0) OR wire_w_man_a_not_zero_w_range142w(0);
	wire_w_lg_w_dataa_range157w159w(0) <= wire_w_dataa_range157w(0) OR wire_w_man_a_not_zero_w_range154w(0);
	wire_w_lg_w_dataa_range163w165w(0) <= wire_w_dataa_range163w(0) OR wire_w_man_a_not_zero_w_range158w(0);
	wire_w_lg_w_dataa_range169w171w(0) <= wire_w_dataa_range169w(0) OR wire_w_man_a_not_zero_w_range164w(0);
	wire_w_lg_w_dataa_range175w177w(0) <= wire_w_dataa_range175w(0) OR wire_w_man_a_not_zero_w_range170w(0);
	wire_w_lg_w_dataa_range181w183w(0) <= wire_w_dataa_range181w(0) OR wire_w_man_a_not_zero_w_range176w(0);
	wire_w_lg_w_dataa_range187w189w(0) <= wire_w_dataa_range187w(0) OR wire_w_man_a_not_zero_w_range182w(0);
	wire_w_lg_w_dataa_range193w195w(0) <= wire_w_dataa_range193w(0) OR wire_w_man_a_not_zero_w_range188w(0);
	wire_w_lg_w_dataa_range87w89w(0) <= wire_w_dataa_range87w(0) OR wire_w_man_a_not_zero_w_range82w(0);
	wire_w_lg_w_dataa_range199w201w(0) <= wire_w_dataa_range199w(0) OR wire_w_man_a_not_zero_w_range194w(0);
	wire_w_lg_w_dataa_range205w207w(0) <= wire_w_dataa_range205w(0) OR wire_w_man_a_not_zero_w_range200w(0);
	wire_w_lg_w_dataa_range211w213w(0) <= wire_w_dataa_range211w(0) OR wire_w_man_a_not_zero_w_range206w(0);
	wire_w_lg_w_dataa_range11w13w(0) <= wire_w_dataa_range11w(0) OR wire_w_exp_a_not_zero_w_range2w(0);
	wire_w_lg_w_dataa_range21w23w(0) <= wire_w_dataa_range21w(0) OR wire_w_exp_a_not_zero_w_range12w(0);
	wire_w_lg_w_dataa_range31w33w(0) <= wire_w_dataa_range31w(0) OR wire_w_exp_a_not_zero_w_range22w(0);
	wire_w_lg_w_dataa_range41w43w(0) <= wire_w_dataa_range41w(0) OR wire_w_exp_a_not_zero_w_range32w(0);
	wire_w_lg_w_dataa_range51w53w(0) <= wire_w_dataa_range51w(0) OR wire_w_exp_a_not_zero_w_range42w(0);
	wire_w_lg_w_dataa_range61w63w(0) <= wire_w_dataa_range61w(0) OR wire_w_exp_a_not_zero_w_range52w(0);
	wire_w_lg_w_dataa_range93w95w(0) <= wire_w_dataa_range93w(0) OR wire_w_man_a_not_zero_w_range88w(0);
	wire_w_lg_w_dataa_range71w73w(0) <= wire_w_dataa_range71w(0) OR wire_w_exp_a_not_zero_w_range62w(0);
	wire_w_lg_w_dataa_range99w101w(0) <= wire_w_dataa_range99w(0) OR wire_w_man_a_not_zero_w_range94w(0);
	wire_w_lg_w_dataa_range105w107w(0) <= wire_w_dataa_range105w(0) OR wire_w_man_a_not_zero_w_range100w(0);
	wire_w_lg_w_dataa_range111w113w(0) <= wire_w_dataa_range111w(0) OR wire_w_man_a_not_zero_w_range106w(0);
	wire_w_lg_w_dataa_range117w119w(0) <= wire_w_dataa_range117w(0) OR wire_w_man_a_not_zero_w_range112w(0);
	wire_w_lg_w_dataa_range123w125w(0) <= wire_w_dataa_range123w(0) OR wire_w_man_a_not_zero_w_range118w(0);
	wire_w_lg_w_dataa_range129w131w(0) <= wire_w_dataa_range129w(0) OR wire_w_man_a_not_zero_w_range124w(0);
	wire_w_lg_w_dataa_range135w137w(0) <= wire_w_dataa_range135w(0) OR wire_w_man_a_not_zero_w_range130w(0);
	wire_w_lg_w_datab_range144w146w(0) <= wire_w_datab_range144w(0) OR wire_w_man_b_not_zero_w_range139w(0);
	wire_w_lg_w_datab_range150w152w(0) <= wire_w_datab_range150w(0) OR wire_w_man_b_not_zero_w_range145w(0);
	wire_w_lg_w_datab_range160w162w(0) <= wire_w_datab_range160w(0) OR wire_w_man_b_not_zero_w_range156w(0);
	wire_w_lg_w_datab_range166w168w(0) <= wire_w_datab_range166w(0) OR wire_w_man_b_not_zero_w_range161w(0);
	wire_w_lg_w_datab_range172w174w(0) <= wire_w_datab_range172w(0) OR wire_w_man_b_not_zero_w_range167w(0);
	wire_w_lg_w_datab_range178w180w(0) <= wire_w_datab_range178w(0) OR wire_w_man_b_not_zero_w_range173w(0);
	wire_w_lg_w_datab_range184w186w(0) <= wire_w_datab_range184w(0) OR wire_w_man_b_not_zero_w_range179w(0);
	wire_w_lg_w_datab_range190w192w(0) <= wire_w_datab_range190w(0) OR wire_w_man_b_not_zero_w_range185w(0);
	wire_w_lg_w_datab_range196w198w(0) <= wire_w_datab_range196w(0) OR wire_w_man_b_not_zero_w_range191w(0);
	wire_w_lg_w_datab_range90w92w(0) <= wire_w_datab_range90w(0) OR wire_w_man_b_not_zero_w_range85w(0);
	wire_w_lg_w_datab_range202w204w(0) <= wire_w_datab_range202w(0) OR wire_w_man_b_not_zero_w_range197w(0);
	wire_w_lg_w_datab_range208w210w(0) <= wire_w_datab_range208w(0) OR wire_w_man_b_not_zero_w_range203w(0);
	wire_w_lg_w_datab_range214w216w(0) <= wire_w_datab_range214w(0) OR wire_w_man_b_not_zero_w_range209w(0);
	wire_w_lg_w_datab_range14w16w(0) <= wire_w_datab_range14w(0) OR wire_w_exp_b_not_zero_w_range5w(0);
	wire_w_lg_w_datab_range24w26w(0) <= wire_w_datab_range24w(0) OR wire_w_exp_b_not_zero_w_range15w(0);
	wire_w_lg_w_datab_range34w36w(0) <= wire_w_datab_range34w(0) OR wire_w_exp_b_not_zero_w_range25w(0);
	wire_w_lg_w_datab_range44w46w(0) <= wire_w_datab_range44w(0) OR wire_w_exp_b_not_zero_w_range35w(0);
	wire_w_lg_w_datab_range54w56w(0) <= wire_w_datab_range54w(0) OR wire_w_exp_b_not_zero_w_range45w(0);
	wire_w_lg_w_datab_range64w66w(0) <= wire_w_datab_range64w(0) OR wire_w_exp_b_not_zero_w_range55w(0);
	wire_w_lg_w_datab_range96w98w(0) <= wire_w_datab_range96w(0) OR wire_w_man_b_not_zero_w_range91w(0);
	wire_w_lg_w_datab_range74w76w(0) <= wire_w_datab_range74w(0) OR wire_w_exp_b_not_zero_w_range65w(0);
	wire_w_lg_w_datab_range102w104w(0) <= wire_w_datab_range102w(0) OR wire_w_man_b_not_zero_w_range97w(0);
	wire_w_lg_w_datab_range108w110w(0) <= wire_w_datab_range108w(0) OR wire_w_man_b_not_zero_w_range103w(0);
	wire_w_lg_w_datab_range114w116w(0) <= wire_w_datab_range114w(0) OR wire_w_man_b_not_zero_w_range109w(0);
	wire_w_lg_w_datab_range120w122w(0) <= wire_w_datab_range120w(0) OR wire_w_man_b_not_zero_w_range115w(0);
	wire_w_lg_w_datab_range126w128w(0) <= wire_w_datab_range126w(0) OR wire_w_man_b_not_zero_w_range121w(0);
	wire_w_lg_w_datab_range132w134w(0) <= wire_w_datab_range132w(0) OR wire_w_man_b_not_zero_w_range127w(0);
	wire_w_lg_w_datab_range138w140w(0) <= wire_w_datab_range138w(0) OR wire_w_man_b_not_zero_w_range133w(0);
	wire_w_lg_w_exp_agb_tmp_w_range265w268w(0) <= wire_w_exp_agb_tmp_w_range265w(0) OR wire_w_exp_eq_gt_grp_range259w(0);
	wire_w_lg_w_exp_agb_tmp_w_range267w270w(0) <= wire_w_exp_agb_tmp_w_range267w(0) OR wire_w_exp_eq_gt_grp_range261w(0);
	wire_w_lg_w_exp_agb_tmp_w_range269w272w(0) <= wire_w_exp_agb_tmp_w_range269w(0) OR wire_w_exp_eq_gt_grp_range263w(0);
	wire_w_lg_w_man_a_not_zero_dffe1_wo_range285w287w(0) <= wire_w_man_a_not_zero_dffe1_wo_range285w(0) OR wire_w_man_a_not_zero_merge_w_range280w(0);
	wire_w_lg_w_man_b_not_zero_dffe1_wo_range288w290w(0) <= wire_w_man_b_not_zero_dffe1_wo_range288w(0) OR wire_w_man_b_not_zero_merge_w_range283w(0);
	wire_w_lg_aligned_dataa_sign_adjusted_dffe2_wo303w(0) <= aligned_dataa_sign_adjusted_dffe2_wo XOR aligned_datab_sign_adjusted_dffe2_wo;
	aclr <= '0';
	alb <= out_alb_dffe3_wo;
	aligned_dataa_sign_adjusted_dffe2_wi <= aligned_dataa_sign_adjusted_w;
	aligned_dataa_sign_adjusted_dffe2_wo <= aligned_dataa_sign_adjusted_dffe2_wi;
	aligned_dataa_sign_adjusted_w <= (aligned_dataa_sign_dffe1_wo AND wire_w_lg_input_dataa_zero_w296w(0));
	aligned_dataa_sign_dffe1_wi <= aligned_dataa_sign_w;
	aligned_dataa_sign_dffe1_wo <= aligned_dataa_sign_dffe1_wi;
	aligned_dataa_sign_w <= dataa(31);
	aligned_dataa_w <= ( dataa(30 DOWNTO 0));
	aligned_datab_sign_adjusted_dffe2_wi <= aligned_datab_sign_adjusted_w;
	aligned_datab_sign_adjusted_dffe2_wo <= aligned_datab_sign_adjusted_dffe2_wi;
	aligned_datab_sign_adjusted_w <= (aligned_datab_sign_dffe1_wo AND wire_w_lg_input_datab_zero_w298w(0));
	aligned_datab_sign_dffe1_wi <= aligned_datab_sign_w;
	aligned_datab_sign_dffe1_wo <= aligned_datab_sign_dffe1_wi;
	aligned_datab_sign_w <= datab(31);
	aligned_datab_w <= ( datab(30 DOWNTO 0));
	both_inputs_zero <= (input_dataa_zero_w AND input_datab_zero_w);
	both_inputs_zero_dffe2_wi <= both_inputs_zero;
	both_inputs_zero_dffe2_wo <= both_inputs_zero_dffe2_wi;
	exp_a_all_one_dffe1_wi <= exp_a_all_one_w(7);
	exp_a_all_one_dffe1_wo <= exp_a_all_one_dffe1_wi;
	exp_a_all_one_w <= ( wire_w_lg_w_dataa_range71w78w & wire_w_lg_w_dataa_range61w68w & wire_w_lg_w_dataa_range51w58w & wire_w_lg_w_dataa_range41w48w & wire_w_lg_w_dataa_range31w38w & wire_w_lg_w_dataa_range21w28w & wire_w_lg_w_dataa_range11w18w & dataa(23));
	exp_a_not_zero_dffe1_wi <= exp_a_not_zero_w(7);
	exp_a_not_zero_dffe1_wo <= exp_a_not_zero_dffe1_wi;
	exp_a_not_zero_w <= ( wire_w_lg_w_dataa_range71w73w & wire_w_lg_w_dataa_range61w63w & wire_w_lg_w_dataa_range51w53w & wire_w_lg_w_dataa_range41w43w & wire_w_lg_w_dataa_range31w33w & wire_w_lg_w_dataa_range21w23w & wire_w_lg_w_dataa_range11w13w & dataa(23));
	exp_aeb <= ( wire_cmpr4_aeb & wire_cmpr3_aeb & wire_cmpr2_aeb & wire_cmpr1_aeb);
	exp_aeb_tmp_w <= ( wire_w_lg_w_exp_aeb_range241w250w & wire_w_lg_w_exp_aeb_range237w248w & wire_w_lg_w_exp_aeb_range233w246w & exp_aeb(0));
	exp_aeb_w <= exp_aeb_tmp_w(3);
	exp_aeb_w_dffe2_wi <= exp_aeb_w;
	exp_aeb_w_dffe2_wo <= exp_aeb_w_dffe2_wi;
	exp_agb <= ( wire_cmpr4_agb & wire_cmpr3_agb & wire_cmpr2_agb & wire_cmpr1_agb);
	exp_agb_tmp_w <= ( wire_w_lg_w_exp_agb_tmp_w_range269w272w & wire_w_lg_w_exp_agb_tmp_w_range267w270w & wire_w_lg_w_exp_agb_tmp_w_range265w268w & exp_eq_gt_grp(0));
	exp_agb_w <= exp_agb_tmp_w(3);
	exp_agb_w_dffe2_wi <= exp_agb_w;
	exp_agb_w_dffe2_wo <= exp_agb_w_dffe2_wi;
	exp_b_all_one_dffe1_wi <= exp_b_all_one_w(7);
	exp_b_all_one_dffe1_wo <= exp_b_all_one_dffe1_wi;
	exp_b_all_one_w <= ( wire_w_lg_w_datab_range74w80w & wire_w_lg_w_datab_range64w70w & wire_w_lg_w_datab_range54w60w & wire_w_lg_w_datab_range44w50w & wire_w_lg_w_datab_range34w40w & wire_w_lg_w_datab_range24w30w & wire_w_lg_w_datab_range14w20w & datab(23));
	exp_b_not_zero_dffe1_wi <= exp_b_not_zero_w(7);
	exp_b_not_zero_dffe1_wo <= exp_b_not_zero_dffe1_wi;
	exp_b_not_zero_w <= ( wire_w_lg_w_datab_range74w76w & wire_w_lg_w_datab_range64w66w & wire_w_lg_w_datab_range54w56w & wire_w_lg_w_datab_range44w46w & wire_w_lg_w_datab_range34w36w & wire_w_lg_w_datab_range24w26w & wire_w_lg_w_datab_range14w16w & datab(23));
	exp_eq_grp <= ( wire_w_lg_w_exp_eq_grp_range253w256w & wire_w_lg_w_exp_eq_grp_range251w254w & exp_aeb(0));
	exp_eq_gt_grp <= ( wire_w_lg_w_exp_eq_grp_range255w264w & wire_w_lg_w_exp_eq_grp_range253w262w & wire_w_lg_w_exp_eq_grp_range251w260w & exp_agb(0));
	flip_outputs_dffe2_wi <= flip_outputs_w;
	flip_outputs_dffe2_wo <= flip_outputs_dffe2_wi;
	flip_outputs_w <= (aligned_dataa_sign_adjusted_w AND aligned_datab_sign_adjusted_w);
	input_dataa_nan_dffe2_wi <= input_dataa_nan_w;
	input_dataa_nan_dffe2_wo <= input_dataa_nan_dffe2_wi;
	input_dataa_nan_w <= (exp_a_all_one_dffe1_wo AND man_a_not_zero_merge_w(1));
	input_dataa_zero_w <= wire_w_lg_exp_a_not_zero_dffe1_wo293w(0);
	input_datab_nan_dffe2_wi <= input_datab_nan_w;
	input_datab_nan_dffe2_wo <= input_datab_nan_dffe2_wi;
	input_datab_nan_w <= (exp_b_all_one_dffe1_wo AND man_b_not_zero_merge_w(1));
	input_datab_zero_w <= wire_w_lg_exp_b_not_zero_dffe1_wo294w(0);
	man_a_not_zero_dffe1_wi <= ( man_a_not_zero_w(22) & man_a_not_zero_w(11));
	man_a_not_zero_dffe1_wo <= man_a_not_zero_dffe1_wi;
	man_a_not_zero_merge_w <= ( wire_w_lg_w_man_a_not_zero_dffe1_wo_range285w287w & man_a_not_zero_dffe1_wo(0));
	man_a_not_zero_w <= ( wire_w_lg_w_dataa_range211w213w & wire_w_lg_w_dataa_range205w207w & wire_w_lg_w_dataa_range199w201w & wire_w_lg_w_dataa_range193w195w & wire_w_lg_w_dataa_range187w189w & wire_w_lg_w_dataa_range181w183w & wire_w_lg_w_dataa_range175w177w & wire_w_lg_w_dataa_range169w171w & wire_w_lg_w_dataa_range163w165w & wire_w_lg_w_dataa_range157w159w & dataa(12) & wire_w_lg_w_dataa_range147w149w & wire_w_lg_w_dataa_range141w143w & wire_w_lg_w_dataa_range135w137w & wire_w_lg_w_dataa_range129w131w & wire_w_lg_w_dataa_range123w125w & wire_w_lg_w_dataa_range117w119w & wire_w_lg_w_dataa_range111w113w & wire_w_lg_w_dataa_range105w107w & wire_w_lg_w_dataa_range99w101w & wire_w_lg_w_dataa_range93w95w & wire_w_lg_w_dataa_range87w89w & dataa(0));
	man_b_not_zero_dffe1_wi <= ( man_b_not_zero_w(22) & man_b_not_zero_w(11));
	man_b_not_zero_dffe1_wo <= man_b_not_zero_dffe1_wi;
	man_b_not_zero_merge_w <= ( wire_w_lg_w_man_b_not_zero_dffe1_wo_range288w290w & man_b_not_zero_dffe1_wo(0));
	man_b_not_zero_w <= ( wire_w_lg_w_datab_range214w216w & wire_w_lg_w_datab_range208w210w & wire_w_lg_w_datab_range202w204w & wire_w_lg_w_datab_range196w198w & wire_w_lg_w_datab_range190w192w & wire_w_lg_w_datab_range184w186w & wire_w_lg_w_datab_range178w180w & wire_w_lg_w_datab_range172w174w & wire_w_lg_w_datab_range166w168w & wire_w_lg_w_datab_range160w162w & datab(12) & wire_w_lg_w_datab_range150w152w & wire_w_lg_w_datab_range144w146w & wire_w_lg_w_datab_range138w140w & wire_w_lg_w_datab_range132w134w & wire_w_lg_w_datab_range126w128w & wire_w_lg_w_datab_range120w122w & wire_w_lg_w_datab_range114w116w & wire_w_lg_w_datab_range108w110w & wire_w_lg_w_datab_range102w104w & wire_w_lg_w_datab_range96w98w & wire_w_lg_w_datab_range90w92w & datab(0));
	out_aeb_w <= (wire_w_lg_w_lg_w304w305w306w(0) AND wire_w_lg_out_unordered_w302w(0));
	out_agb_w <= (((wire_w316w(0) OR (wire_w_lg_exp_agb_w_dffe2_wo314w(0) AND wire_w_lg_both_inputs_zero_dffe2_wo312w(0))) OR (wire_w_lg_flip_outputs_dffe2_wo310w(0) AND wire_w_lg_out_aeb_w308w(0))) AND wire_w_lg_out_unordered_w302w(0));
	out_alb_dffe3_wi <= out_alb_w;
	out_alb_dffe3_wo <= out_alb_w_dffe3;
	out_alb_w <= ((wire_w_lg_out_agb_w320w(0) AND wire_w_lg_out_aeb_w308w(0)) AND wire_w_lg_out_unordered_w302w(0));
	out_unordered_w <= (input_dataa_nan_dffe2_wo OR input_datab_nan_dffe2_wo);
	wire_w_dataa_range141w(0) <= dataa(10);
	wire_w_dataa_range147w(0) <= dataa(11);
	wire_w_dataa_range157w(0) <= dataa(13);
	wire_w_dataa_range163w(0) <= dataa(14);
	wire_w_dataa_range169w(0) <= dataa(15);
	wire_w_dataa_range175w(0) <= dataa(16);
	wire_w_dataa_range181w(0) <= dataa(17);
	wire_w_dataa_range187w(0) <= dataa(18);
	wire_w_dataa_range193w(0) <= dataa(19);
	wire_w_dataa_range87w(0) <= dataa(1);
	wire_w_dataa_range199w(0) <= dataa(20);
	wire_w_dataa_range205w(0) <= dataa(21);
	wire_w_dataa_range211w(0) <= dataa(22);
	wire_w_dataa_range11w(0) <= dataa(24);
	wire_w_dataa_range21w(0) <= dataa(25);
	wire_w_dataa_range31w(0) <= dataa(26);
	wire_w_dataa_range41w(0) <= dataa(27);
	wire_w_dataa_range51w(0) <= dataa(28);
	wire_w_dataa_range61w(0) <= dataa(29);
	wire_w_dataa_range93w(0) <= dataa(2);
	wire_w_dataa_range71w(0) <= dataa(30);
	wire_w_dataa_range99w(0) <= dataa(3);
	wire_w_dataa_range105w(0) <= dataa(4);
	wire_w_dataa_range111w(0) <= dataa(5);
	wire_w_dataa_range117w(0) <= dataa(6);
	wire_w_dataa_range123w(0) <= dataa(7);
	wire_w_dataa_range129w(0) <= dataa(8);
	wire_w_dataa_range135w(0) <= dataa(9);
	wire_w_datab_range144w(0) <= datab(10);
	wire_w_datab_range150w(0) <= datab(11);
	wire_w_datab_range160w(0) <= datab(13);
	wire_w_datab_range166w(0) <= datab(14);
	wire_w_datab_range172w(0) <= datab(15);
	wire_w_datab_range178w(0) <= datab(16);
	wire_w_datab_range184w(0) <= datab(17);
	wire_w_datab_range190w(0) <= datab(18);
	wire_w_datab_range196w(0) <= datab(19);
	wire_w_datab_range90w(0) <= datab(1);
	wire_w_datab_range202w(0) <= datab(20);
	wire_w_datab_range208w(0) <= datab(21);
	wire_w_datab_range214w(0) <= datab(22);
	wire_w_datab_range14w(0) <= datab(24);
	wire_w_datab_range24w(0) <= datab(25);
	wire_w_datab_range34w(0) <= datab(26);
	wire_w_datab_range44w(0) <= datab(27);
	wire_w_datab_range54w(0) <= datab(28);
	wire_w_datab_range64w(0) <= datab(29);
	wire_w_datab_range96w(0) <= datab(2);
	wire_w_datab_range74w(0) <= datab(30);
	wire_w_datab_range102w(0) <= datab(3);
	wire_w_datab_range108w(0) <= datab(4);
	wire_w_datab_range114w(0) <= datab(5);
	wire_w_datab_range120w(0) <= datab(6);
	wire_w_datab_range126w(0) <= datab(7);
	wire_w_datab_range132w(0) <= datab(8);
	wire_w_datab_range138w(0) <= datab(9);
	wire_w_exp_a_all_one_w_range7w(0) <= exp_a_all_one_w(0);
	wire_w_exp_a_all_one_w_range17w(0) <= exp_a_all_one_w(1);
	wire_w_exp_a_all_one_w_range27w(0) <= exp_a_all_one_w(2);
	wire_w_exp_a_all_one_w_range37w(0) <= exp_a_all_one_w(3);
	wire_w_exp_a_all_one_w_range47w(0) <= exp_a_all_one_w(4);
	wire_w_exp_a_all_one_w_range57w(0) <= exp_a_all_one_w(5);
	wire_w_exp_a_all_one_w_range67w(0) <= exp_a_all_one_w(6);
	wire_w_exp_a_not_zero_w_range2w(0) <= exp_a_not_zero_w(0);
	wire_w_exp_a_not_zero_w_range12w(0) <= exp_a_not_zero_w(1);
	wire_w_exp_a_not_zero_w_range22w(0) <= exp_a_not_zero_w(2);
	wire_w_exp_a_not_zero_w_range32w(0) <= exp_a_not_zero_w(3);
	wire_w_exp_a_not_zero_w_range42w(0) <= exp_a_not_zero_w(4);
	wire_w_exp_a_not_zero_w_range52w(0) <= exp_a_not_zero_w(5);
	wire_w_exp_a_not_zero_w_range62w(0) <= exp_a_not_zero_w(6);
	wire_w_exp_aeb_range233w(0) <= exp_aeb(1);
	wire_w_exp_aeb_range237w(0) <= exp_aeb(2);
	wire_w_exp_aeb_range241w(0) <= exp_aeb(3);
	wire_w_exp_aeb_tmp_w_range243w(0) <= exp_aeb_tmp_w(0);
	wire_w_exp_aeb_tmp_w_range245w(0) <= exp_aeb_tmp_w(1);
	wire_w_exp_aeb_tmp_w_range247w(0) <= exp_aeb_tmp_w(2);
	wire_w_exp_agb_range234w(0) <= exp_agb(1);
	wire_w_exp_agb_range238w(0) <= exp_agb(2);
	wire_w_exp_agb_range242w(0) <= exp_agb(3);
	wire_w_exp_agb_tmp_w_range265w(0) <= exp_agb_tmp_w(0);
	wire_w_exp_agb_tmp_w_range267w(0) <= exp_agb_tmp_w(1);
	wire_w_exp_agb_tmp_w_range269w(0) <= exp_agb_tmp_w(2);
	wire_w_exp_b_all_one_w_range9w(0) <= exp_b_all_one_w(0);
	wire_w_exp_b_all_one_w_range19w(0) <= exp_b_all_one_w(1);
	wire_w_exp_b_all_one_w_range29w(0) <= exp_b_all_one_w(2);
	wire_w_exp_b_all_one_w_range39w(0) <= exp_b_all_one_w(3);
	wire_w_exp_b_all_one_w_range49w(0) <= exp_b_all_one_w(4);
	wire_w_exp_b_all_one_w_range59w(0) <= exp_b_all_one_w(5);
	wire_w_exp_b_all_one_w_range69w(0) <= exp_b_all_one_w(6);
	wire_w_exp_b_not_zero_w_range5w(0) <= exp_b_not_zero_w(0);
	wire_w_exp_b_not_zero_w_range15w(0) <= exp_b_not_zero_w(1);
	wire_w_exp_b_not_zero_w_range25w(0) <= exp_b_not_zero_w(2);
	wire_w_exp_b_not_zero_w_range35w(0) <= exp_b_not_zero_w(3);
	wire_w_exp_b_not_zero_w_range45w(0) <= exp_b_not_zero_w(4);
	wire_w_exp_b_not_zero_w_range55w(0) <= exp_b_not_zero_w(5);
	wire_w_exp_b_not_zero_w_range65w(0) <= exp_b_not_zero_w(6);
	wire_w_exp_eq_grp_range251w(0) <= exp_eq_grp(0);
	wire_w_exp_eq_grp_range253w(0) <= exp_eq_grp(1);
	wire_w_exp_eq_grp_range255w(0) <= exp_eq_grp(2);
	wire_w_exp_eq_gt_grp_range259w(0) <= exp_eq_gt_grp(1);
	wire_w_exp_eq_gt_grp_range261w(0) <= exp_eq_gt_grp(2);
	wire_w_exp_eq_gt_grp_range263w(0) <= exp_eq_gt_grp(3);
	wire_w_man_a_not_zero_dffe1_wo_range285w(0) <= man_a_not_zero_dffe1_wo(1);
	wire_w_man_a_not_zero_merge_w_range280w(0) <= man_a_not_zero_merge_w(0);
	wire_w_man_a_not_zero_w_range82w(0) <= man_a_not_zero_w(0);
	wire_w_man_a_not_zero_w_range142w(0) <= man_a_not_zero_w(10);
	wire_w_man_a_not_zero_w_range154w(0) <= man_a_not_zero_w(12);
	wire_w_man_a_not_zero_w_range158w(0) <= man_a_not_zero_w(13);
	wire_w_man_a_not_zero_w_range164w(0) <= man_a_not_zero_w(14);
	wire_w_man_a_not_zero_w_range170w(0) <= man_a_not_zero_w(15);
	wire_w_man_a_not_zero_w_range176w(0) <= man_a_not_zero_w(16);
	wire_w_man_a_not_zero_w_range182w(0) <= man_a_not_zero_w(17);
	wire_w_man_a_not_zero_w_range188w(0) <= man_a_not_zero_w(18);
	wire_w_man_a_not_zero_w_range194w(0) <= man_a_not_zero_w(19);
	wire_w_man_a_not_zero_w_range88w(0) <= man_a_not_zero_w(1);
	wire_w_man_a_not_zero_w_range200w(0) <= man_a_not_zero_w(20);
	wire_w_man_a_not_zero_w_range206w(0) <= man_a_not_zero_w(21);
	wire_w_man_a_not_zero_w_range94w(0) <= man_a_not_zero_w(2);
	wire_w_man_a_not_zero_w_range100w(0) <= man_a_not_zero_w(3);
	wire_w_man_a_not_zero_w_range106w(0) <= man_a_not_zero_w(4);
	wire_w_man_a_not_zero_w_range112w(0) <= man_a_not_zero_w(5);
	wire_w_man_a_not_zero_w_range118w(0) <= man_a_not_zero_w(6);
	wire_w_man_a_not_zero_w_range124w(0) <= man_a_not_zero_w(7);
	wire_w_man_a_not_zero_w_range130w(0) <= man_a_not_zero_w(8);
	wire_w_man_a_not_zero_w_range136w(0) <= man_a_not_zero_w(9);
	wire_w_man_b_not_zero_dffe1_wo_range288w(0) <= man_b_not_zero_dffe1_wo(1);
	wire_w_man_b_not_zero_merge_w_range283w(0) <= man_b_not_zero_merge_w(0);
	wire_w_man_b_not_zero_w_range85w(0) <= man_b_not_zero_w(0);
	wire_w_man_b_not_zero_w_range145w(0) <= man_b_not_zero_w(10);
	wire_w_man_b_not_zero_w_range156w(0) <= man_b_not_zero_w(12);
	wire_w_man_b_not_zero_w_range161w(0) <= man_b_not_zero_w(13);
	wire_w_man_b_not_zero_w_range167w(0) <= man_b_not_zero_w(14);
	wire_w_man_b_not_zero_w_range173w(0) <= man_b_not_zero_w(15);
	wire_w_man_b_not_zero_w_range179w(0) <= man_b_not_zero_w(16);
	wire_w_man_b_not_zero_w_range185w(0) <= man_b_not_zero_w(17);
	wire_w_man_b_not_zero_w_range191w(0) <= man_b_not_zero_w(18);
	wire_w_man_b_not_zero_w_range197w(0) <= man_b_not_zero_w(19);
	wire_w_man_b_not_zero_w_range91w(0) <= man_b_not_zero_w(1);
	wire_w_man_b_not_zero_w_range203w(0) <= man_b_not_zero_w(20);
	wire_w_man_b_not_zero_w_range209w(0) <= man_b_not_zero_w(21);
	wire_w_man_b_not_zero_w_range97w(0) <= man_b_not_zero_w(2);
	wire_w_man_b_not_zero_w_range103w(0) <= man_b_not_zero_w(3);
	wire_w_man_b_not_zero_w_range109w(0) <= man_b_not_zero_w(4);
	wire_w_man_b_not_zero_w_range115w(0) <= man_b_not_zero_w(5);
	wire_w_man_b_not_zero_w_range121w(0) <= man_b_not_zero_w(6);
	wire_w_man_b_not_zero_w_range127w(0) <= man_b_not_zero_w(7);
	wire_w_man_b_not_zero_w_range133w(0) <= man_b_not_zero_w(8);
	wire_w_man_b_not_zero_w_range139w(0) <= man_b_not_zero_w(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN out_alb_w_dffe3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN out_alb_w_dffe3 <= out_alb_dffe3_wi;
			END IF;
		END IF;
	END PROCESS;
	cmpr1 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr1_aeb,
		agb => wire_cmpr1_agb,
		dataa => aligned_dataa_w(30 DOWNTO 23),
		datab => aligned_datab_w(30 DOWNTO 23)
	  );
	cmpr2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr2_aeb,
		agb => wire_cmpr2_agb,
		dataa => aligned_dataa_w(22 DOWNTO 15),
		datab => aligned_datab_w(22 DOWNTO 15)
	  );
	cmpr3 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aeb => wire_cmpr3_aeb,
		agb => wire_cmpr3_agb,
		dataa => aligned_dataa_w(14 DOWNTO 7),
		datab => aligned_datab_w(14 DOWNTO 7)
	  );
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 7
	  )
	  PORT MAP ( 
		aeb => wire_cmpr4_aeb,
		agb => wire_cmpr4_agb,
		dataa => aligned_dataa_w(6 DOWNTO 0),
		datab => aligned_datab_w(6 DOWNTO 0)
	  );

 END RTL; --CompareALessB_altfp_compare_ksb
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CompareALessB IS
	PORT
	(
		clk_en		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		alb		: OUT STD_LOGIC 
	);
END CompareALessB;


ARCHITECTURE RTL OF comparealessb IS

	SIGNAL sub_wire0	: STD_LOGIC ;



	COMPONENT CompareALessB_altfp_compare_ksb
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			alb	: OUT STD_LOGIC ;
			clk_en	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	alb    <= sub_wire0;

	CompareALessB_altfp_compare_ksb_component : CompareALessB_altfp_compare_ksb
	PORT MAP (
		dataa => dataa,
		datab => datab,
		clk_en => clk_en,
		clock => clock,
		alb => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: alb 0 0 0 0 OUTPUT NODEFVAL "alb"
-- Retrieval info: USED_PORT: clk_en 0 0 0 0 INPUT NODEFVAL "clk_en"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL "datab[31..0]"
-- Retrieval info: CONNECT: @clk_en 0 0 0 0 clk_en 0 0 0 0
-- Retrieval info: CONNECT: alb 0 0 0 0 @alb 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL CompareALessB.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CompareALessB.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CompareALessB.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CompareALessB.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL CompareALessB_inst.vhd TRUE
-- Retrieval info: LIB_FILE: lpm

