CompareAMenorB_inst : CompareAMenorB PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		alb	 => alb_sig
	);
