-- megafunction wizard: %PARALLEL_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: parallel_add 

-- ============================================================
-- File Name: ParallelAdd.vhd
-- Megafunction Name(s):
-- 			parallel_add
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.1.0 Build 196 10/24/2016 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2016  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Intel and sold by Intel or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY ParallelAdd IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END ParallelAdd;


ARCHITECTURE SYN OF paralleladd IS

--	type ALTERA_MF_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: ALTERA_MF_LOGIC_2D (7 DOWNTO 0, 0 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (3 DOWNTO 0);

BEGIN
	sub_wire8    <= data0x(0 DOWNTO 0);
	sub_wire7    <= data1x(0 DOWNTO 0);
	sub_wire6    <= data2x(0 DOWNTO 0);
	sub_wire5    <= data3x(0 DOWNTO 0);
	sub_wire4    <= data4x(0 DOWNTO 0);
	sub_wire3    <= data5x(0 DOWNTO 0);
	sub_wire2    <= data6x(0 DOWNTO 0);
	sub_wire0    <= data7x(0 DOWNTO 0);
	sub_wire1(7, 0)    <= sub_wire0(0);
	sub_wire1(6, 0)    <= sub_wire2(0);
	sub_wire1(5, 0)    <= sub_wire3(0);
	sub_wire1(4, 0)    <= sub_wire4(0);
	sub_wire1(3, 0)    <= sub_wire5(0);
	sub_wire1(2, 0)    <= sub_wire6(0);
	sub_wire1(1, 0)    <= sub_wire7(0);
	sub_wire1(0, 0)    <= sub_wire8(0);
	result    <= sub_wire9(3 DOWNTO 0);

	parallel_add_component : parallel_add
	GENERIC MAP (
		msw_subtract => "NO",
		pipeline => 0,
		representation => "UNSIGNED",
		result_alignment => "LSB",
		shift => 0,
		size => 8,
		width => 1,
		widthr => 4,
		lpm_type => "parallel_add"
	)
	PORT MAP (
		data => sub_wire1,
		result => sub_wire9
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
-- Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
-- Retrieval info: CONSTANT: SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: SIZE NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTHR NUMERIC "4"
-- Retrieval info: USED_PORT: data0x 0 0 1 0 INPUT NODEFVAL "data0x[0..0]"
-- Retrieval info: USED_PORT: data1x 0 0 1 0 INPUT NODEFVAL "data1x[0..0]"
-- Retrieval info: USED_PORT: data2x 0 0 1 0 INPUT NODEFVAL "data2x[0..0]"
-- Retrieval info: USED_PORT: data3x 0 0 1 0 INPUT NODEFVAL "data3x[0..0]"
-- Retrieval info: USED_PORT: data4x 0 0 1 0 INPUT NODEFVAL "data4x[0..0]"
-- Retrieval info: USED_PORT: data5x 0 0 1 0 INPUT NODEFVAL "data5x[0..0]"
-- Retrieval info: USED_PORT: data6x 0 0 1 0 INPUT NODEFVAL "data6x[0..0]"
-- Retrieval info: USED_PORT: data7x 0 0 1 0 INPUT NODEFVAL "data7x[0..0]"
-- Retrieval info: USED_PORT: result 0 0 4 0 OUTPUT NODEFVAL "result[3..0]"
-- Retrieval info: CONNECT: @data 1 0 1 0 data0x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 1 1 0 data1x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 2 1 0 data2x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 3 1 0 data3x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 4 1 0 data4x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 5 1 0 data5x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 6 1 0 data6x 0 0 1 0
-- Retrieval info: CONNECT: @data 1 7 1 0 data7x 0 0 1 0
-- Retrieval info: CONNECT: result 0 0 4 0 @result 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ParallelAdd.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ParallelAdd.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ParallelAdd.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ParallelAdd.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ParallelAdd_inst.vhd TRUE
-- Retrieval info: LIB_FILE: altera_mf
