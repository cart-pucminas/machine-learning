ShiftReg_FP_inst : ShiftReg_FP PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		shiftout	 => shiftout_sig
	);
